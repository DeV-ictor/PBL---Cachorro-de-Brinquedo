module display (
	input clk,
	output reg q
);

	initial begin
	end
	
	always @(posedge clk or negedge clk) begin
		
		
	
	end

endmodule