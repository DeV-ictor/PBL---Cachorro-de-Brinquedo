module t_ff (
  input clk, t, reset,
  output reg q
);

  // Inicialização do valor de q
  initial begin
    q = 0;
  end

  // Lógica do flip-flop T
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q <= 0; // Reinicialização 
    end else begin
      if (t) begin
			q <= 1;
		end
    end
  end

endmodule
